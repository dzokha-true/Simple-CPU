module register(d, clk, en, rst, q);
		input [15:0] d;
		input clk, rst, en;
		output reg [15:0] q;
		
		parameter num_bits = 16;
		
		always @ (posedge clk or posedge rst) begin
			if (rst == 1'b1)
				q_out <= {num_bits{1'b0}};
			else begin
				if (en == 1'b1)
					q <= d;
				else
					q <= q;
			end
		end

endmodule
