module state_reg(d, clk, rst, q);
		input [4:0] d;
		input clk, rst;
		output reg [4:0] q;
		
		parameter num_bits = 5;
		
		always @ (posedge clk or posedge rst) begin
			if (rst == 1'b1)
				q_out <= {num_bits{1'b0}};
			else begin
				if (en == 1'b1)
					q <= d;
				else
					q <= q;
			end
		end

endmodule